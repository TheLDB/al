module compiler

pub struct AST {
	//
}

fn (ast AST) str() string {
	return print(&ast)
}
