module compiler

import math

const (
	single_quote = `'`
	// char used as number separator
	num_sep      = `_`
	b_lf         = 10
	b_cr         = 13
	backslash    = `\\`
)

[minify]
pub struct ScannerState {
pub mut:
	nr_lines                    int // Total number of lines
	last_nl_pos                 int = -1 // Used to calculate column
	tidx                        int
	pos                         int
	line                        int
	should_abort                bool
	is_crlf                     bool
	is_inside_string            bool
	is_string_interpolation_end bool
}

[minify]
pub struct Scanner {
pub:
	absolute_file_path string // The absolute path of the file
	text               string // The whole text of the file
pub mut:
	state      ScannerState
	all_tokens []Token = []Token{}
mut:
	messages []Message = []Message{} // Messages generated by the scanner
}

[inline]
fn (mut s Scanner) new_token(tok_kind Kind, lit string, len int) Token {
	// cidx := s.tidx
	s.state.tidx++

	return Token{
		kind: tok_kind
		lit: lit
		line: s.state.line
		col: math.max(1, s.current_column() - len + 1)
		scanner_pos: s.state.pos - len + 1
		len: len
	}
}

pub fn (mut s Scanner) text_scan() Token {
	for {
		s.state.pos++

		if s.state.is_inside_string {
			s.skip_whitespace()
		}

		if s.state.pos >= s.text.len || s.state.should_abort {
			return s.end_of_file()
		}

		if s.state.is_string_interpolation_end {
			if s.text[s.state.pos] == s.state.quote {
				s.is_inter_end = false
				return s.new_token(.string, '', 1)
			}

			s.state.is_string_interpolation_end = falser
			ident_string := s.ident_string()

			return s.new_token(.string, ident_string, ident_string.len + 2) // + two quotes
		}
	}

	return s.new_token(.eof, '', 1)
}

fn (s &Scanner) current_column() int {
	return s.state.pos - s.state.last_nl_pos
}

pub fn new_scanner(absolute_file_path string, text string) Scanner {
	return Scanner{
		absolute_file_path: absolute_file_path
		text: text
	}
}

pub fn (s &Scanner) peek() byte {
	return s.text[s.state.pos]
}

pub fn (s &Scanner) look_ahead(n int) string {
	return (s.text[s.state.pos..s.state.pos + n]).str()
}

fn (mut s Scanner) end_of_file() Token {
	if s.state.pos != s.text.len {
		s.inc_line_number()
	}

	s.state.pos = s.text.len

	return s.new_eof_token()
}

[inline]
fn (mut s Scanner) inc_line_number() {
	if s.state.is_crlf {
		s.state.last_nl_pos++
	}

	s.state.line++

	if s.state.line > s.state.nr_lines {
		s.state.nr_lines = s.state.line
	}
}

[direct_array_access; inline]
fn (mut s Scanner) skip_whitespace() {
	for s.state.pos < s.text.len {
		c := s.text[s.state.pos]

		// Tabs
		if c == 9 {
			s.state.pos++
			continue
		}

		if !(c == 32 || (c > 8 && c < 14) || (c == 0x85) || (c == 0xa0)) {
			return
		}

		c_is_nl := c == compiler.b_cr || c == compiler.b_lf

		if s.state.pos + 1 < s.text.len && c == compiler.b_cr
			&& s.text[s.state.pos + 1] == compiler.b_lf {
			s.state.is_crlf = true
		}

		// Count \r\n as one line
		if c_is_nl && !(s.state.pos > 0 && s.text[s.state.pos - 1] == compiler.b_cr
			&& c == compiler.b_lf) {
			s.inc_line_number()
		}

		s.state.pos++
	}
}

pub fn (mut s Scanner) scan() {
	for {
		t := s.text_scan()

		s.all_tokens << t

		if t.kind == .eof || s.state.should_abort {
			break
		}
	}
}

[inline]
fn (s &Scanner) new_eof_token() Token {
	return Token{
		kind: .eof
		lit: ''
		line: s.state.line + 1
		col: s.current_column()
		len: 1
	}
}
