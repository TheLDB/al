module compiler

// TODO: Implement this function
pub fn print(ast &AST) string {
	return ''
}
